library verilog;
use verilog.vl_types.all;
entity proj_vlg_vec_tst is
end proj_vlg_vec_tst;
